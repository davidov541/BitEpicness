`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:04:49 02/20/2011 
// Design Name: 
// Module Name:    receiveSD 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module receiveSD(input clock, input reset, input enable, input SDin, output reg [7:0] received, output done);


	reg [1:0] state, nextState;
	wire resetReceived, save;
	
	reg [2:0] count;
	wire countDone;
	
	assign countDone = (count == 3'b000);
	assign resetReceived = (state == 2'b01);
	assign save = (state == 2'b10);
	assign done = (state == 2'b11);
	
	
	always @(posedge clock, posedge reset)
	if (reset)
		begin
			state <= 2'b00;
			received <= 8'b00000000;
			count <= 3'b000;
		end
	else
		begin
			state <= nextState;
			received <= (resetReceived) ? 8'b00000000 : (save) ? {received[6:0], SDin} : received;
			count <= (resetReceived) ? 3'b110 : (countDone) ? 3'b000 : count - 1;
		end
		
	always @(*)
	case(state)
	2'b00: nextState = (enable) ? 2'b01 : 2'b00;
	2'b01: nextState = (SDin == 1'b0) ? 2'b10 : 2'b01;
	2'b10: nextState = (countDone) ? 2'b11 : 2'b10;
	2'b11: nextState = 2'b00;
	default: nextState = 2'b00;
	endcase
	
endmodule
