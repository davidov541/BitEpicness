// Encoder32bit
//
// Encodes a 32 inputs into a 5 bit number
module Encoder32bit(
    input [31:0] dataIn,
    output [4:0] dataOut
    );


	assign dataOut = (dataIn == 32'b00000000000000000000000000000000) ? 5'b00000 :
	(dataIn == 32'b00000000000000000000000000000001) ? 5'b00000 :
	(dataIn == 32'b00000000000000000000000000000010) ? 5'b00001 :
	(dataIn == 32'b00000000000000000000000000000100) ? 5'b00010 :
	(dataIn == 32'b00000000000000000000000000001000) ? 5'b00011 :
	(dataIn == 32'b00000000000000000000000000010000) ? 5'b00100 :
	(dataIn == 32'b00000000000000000000000000100000) ? 5'b00101 :
	(dataIn == 32'b00000000000000000000000001000000) ? 5'b00110 :
	(dataIn == 32'b00000000000000000000000010000000) ? 5'b00111 :
	(dataIn == 32'b00000000000000000000000100000000) ? 5'b01000 :
	(dataIn == 32'b00000000000000000000001000000000) ? 5'b01001 :
	(dataIn == 32'b00000000000000000000010000000000) ? 5'b01010 :
	(dataIn == 32'b00000000000000000000100000000000) ? 5'b01011 :
	(dataIn == 32'b00000000000000000001000000000000) ? 5'b01100 :
	(dataIn == 32'b00000000000000000010000000000000) ? 5'b01101 :
	(dataIn == 32'b00000000000000000100000000000000) ? 5'b01110 :
	(dataIn == 32'b00000000000000001000000000000000) ? 5'b01111 :
	(dataIn == 32'b00000000000000010000000000000000) ? 5'b10000 :
	(dataIn == 32'b00000000000000100000000000000000) ? 5'b10001 :
	(dataIn == 32'b00000000000001000000000000000000) ? 5'b10010 :
	(dataIn == 32'b00000000000010000000000000000000) ? 5'b10011 :
	(dataIn == 32'b00000000000100000000000000000000) ? 5'b10100 :
	(dataIn == 32'b00000000001000000000000000000000) ? 5'b10101 :
	(dataIn == 32'b00000000010000000000000000000000) ? 5'b10110 :
	(dataIn == 32'b00000000100000000000000000000000) ? 5'b10111 :
	(dataIn == 32'b00000001000000000000000000000000) ? 5'b11000 :
	(dataIn == 32'b00000010000000000000000000000000) ? 5'b11001 :
	(dataIn == 32'b00000100000000000000000000000000) ? 5'b11010 :
	(dataIn == 32'b00001000000000000000000000000000) ? 5'b11011 :
	(dataIn == 32'b00010000000000000000000000000000) ? 5'b11100 :
	(dataIn == 32'b00100000000000000000000000000000) ? 5'b11101 :
	(dataIn == 32'b01000000000000000000000000000000) ? 5'b11110 :
	(dataIn == 32'b10000000000000000000000000000000) ? 5'b11111 : 5'bXXXXX;
	
		

endmodule
